VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO arbiterpuf
  CLASS BLOCK ;
  FOREIGN arbiterpuf ;
  ORIGIN 0.000 0.000 ;
  SIZE 400.000 BY 400.000 ;
  PIN ichallenge[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.130 396.000 34.410 400.000 ;
    END
  END ichallenge[0]
  PIN ichallenge[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.930 396.000 255.210 400.000 ;
    END
  END ichallenge[10]
  PIN ichallenge[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.010 396.000 277.290 400.000 ;
    END
  END ichallenge[11]
  PIN ichallenge[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.090 396.000 299.370 400.000 ;
    END
  END ichallenge[12]
  PIN ichallenge[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 321.170 396.000 321.450 400.000 ;
    END
  END ichallenge[13]
  PIN ichallenge[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 343.250 396.000 343.530 400.000 ;
    END
  END ichallenge[14]
  PIN ichallenge[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 365.330 396.000 365.610 400.000 ;
    END
  END ichallenge[15]
  PIN ichallenge[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.210 396.000 56.490 400.000 ;
    END
  END ichallenge[1]
  PIN ichallenge[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.290 396.000 78.570 400.000 ;
    END
  END ichallenge[2]
  PIN ichallenge[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.370 396.000 100.650 400.000 ;
    END
  END ichallenge[3]
  PIN ichallenge[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.450 396.000 122.730 400.000 ;
    END
  END ichallenge[4]
  PIN ichallenge[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.530 396.000 144.810 400.000 ;
    END
  END ichallenge[5]
  PIN ichallenge[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 166.610 396.000 166.890 400.000 ;
    END
  END ichallenge[6]
  PIN ichallenge[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 188.690 396.000 188.970 400.000 ;
    END
  END ichallenge[7]
  PIN ichallenge[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 210.770 396.000 211.050 400.000 ;
    END
  END ichallenge[8]
  PIN ichallenge[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 232.850 396.000 233.130 400.000 ;
    END
  END ichallenge[9]
  PIN ipulse
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.050 396.000 12.330 400.000 ;
    END
  END ipulse
  PIN oresponse
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 387.410 396.000 387.690 400.000 ;
    END
  END oresponse
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 389.200 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 389.200 ;
    END
  END vssd1
  OBS
      LAYER nwell ;
        RECT 5.330 387.545 394.410 389.150 ;
        RECT 5.330 382.105 394.410 384.935 ;
        RECT 5.330 376.665 394.410 379.495 ;
        RECT 5.330 371.225 394.410 374.055 ;
        RECT 5.330 365.785 394.410 368.615 ;
        RECT 5.330 360.345 394.410 363.175 ;
        RECT 5.330 354.905 394.410 357.735 ;
        RECT 5.330 349.465 394.410 352.295 ;
        RECT 5.330 344.025 394.410 346.855 ;
        RECT 5.330 338.585 394.410 341.415 ;
        RECT 5.330 333.145 394.410 335.975 ;
        RECT 5.330 327.705 394.410 330.535 ;
        RECT 5.330 322.265 394.410 325.095 ;
        RECT 5.330 316.825 394.410 319.655 ;
        RECT 5.330 311.385 394.410 314.215 ;
        RECT 5.330 305.945 394.410 308.775 ;
        RECT 5.330 300.505 394.410 303.335 ;
        RECT 5.330 295.065 394.410 297.895 ;
        RECT 5.330 289.625 394.410 292.455 ;
        RECT 5.330 284.185 394.410 287.015 ;
        RECT 5.330 278.745 394.410 281.575 ;
        RECT 5.330 273.305 394.410 276.135 ;
        RECT 5.330 267.865 394.410 270.695 ;
        RECT 5.330 262.425 394.410 265.255 ;
        RECT 5.330 256.985 394.410 259.815 ;
        RECT 5.330 251.545 394.410 254.375 ;
        RECT 5.330 246.105 394.410 248.935 ;
        RECT 5.330 240.665 394.410 243.495 ;
        RECT 5.330 235.225 394.410 238.055 ;
        RECT 5.330 229.785 394.410 232.615 ;
        RECT 5.330 224.345 394.410 227.175 ;
        RECT 5.330 218.905 394.410 221.735 ;
        RECT 5.330 213.465 394.410 216.295 ;
        RECT 5.330 208.025 394.410 210.855 ;
        RECT 5.330 202.585 394.410 205.415 ;
        RECT 5.330 197.145 394.410 199.975 ;
        RECT 5.330 191.705 394.410 194.535 ;
        RECT 5.330 186.265 394.410 189.095 ;
        RECT 5.330 180.825 394.410 183.655 ;
        RECT 5.330 175.385 394.410 178.215 ;
        RECT 5.330 169.945 394.410 172.775 ;
        RECT 5.330 164.505 394.410 167.335 ;
        RECT 5.330 159.065 394.410 161.895 ;
        RECT 5.330 153.625 394.410 156.455 ;
        RECT 5.330 148.185 394.410 151.015 ;
        RECT 5.330 142.745 394.410 145.575 ;
        RECT 5.330 137.305 394.410 140.135 ;
        RECT 5.330 131.865 394.410 134.695 ;
        RECT 5.330 126.425 394.410 129.255 ;
        RECT 5.330 120.985 394.410 123.815 ;
        RECT 5.330 115.545 394.410 118.375 ;
        RECT 5.330 110.105 394.410 112.935 ;
        RECT 5.330 104.665 394.410 107.495 ;
        RECT 5.330 99.225 394.410 102.055 ;
        RECT 5.330 93.785 394.410 96.615 ;
        RECT 5.330 88.345 394.410 91.175 ;
        RECT 5.330 82.905 394.410 85.735 ;
        RECT 5.330 77.465 394.410 80.295 ;
        RECT 5.330 72.025 394.410 74.855 ;
        RECT 5.330 66.585 394.410 69.415 ;
        RECT 5.330 61.145 394.410 63.975 ;
        RECT 5.330 55.705 394.410 58.535 ;
        RECT 5.330 50.265 394.410 53.095 ;
        RECT 5.330 44.825 394.410 47.655 ;
        RECT 5.330 39.385 394.410 42.215 ;
        RECT 5.330 33.945 394.410 36.775 ;
        RECT 5.330 28.505 394.410 31.335 ;
        RECT 5.330 23.065 394.410 25.895 ;
        RECT 5.330 17.625 394.410 20.455 ;
        RECT 5.330 12.185 394.410 15.015 ;
      LAYER li1 ;
        RECT 5.520 10.795 394.220 389.045 ;
      LAYER met1 ;
        RECT 5.520 10.640 394.220 389.200 ;
      LAYER met2 ;
        RECT 12.610 395.720 33.850 396.000 ;
        RECT 34.690 395.720 55.930 396.000 ;
        RECT 56.770 395.720 78.010 396.000 ;
        RECT 78.850 395.720 100.090 396.000 ;
        RECT 100.930 395.720 122.170 396.000 ;
        RECT 123.010 395.720 144.250 396.000 ;
        RECT 145.090 395.720 166.330 396.000 ;
        RECT 167.170 395.720 188.410 396.000 ;
        RECT 189.250 395.720 210.490 396.000 ;
        RECT 211.330 395.720 232.570 396.000 ;
        RECT 233.410 395.720 254.650 396.000 ;
        RECT 255.490 395.720 276.730 396.000 ;
        RECT 277.570 395.720 298.810 396.000 ;
        RECT 299.650 395.720 320.890 396.000 ;
        RECT 321.730 395.720 342.970 396.000 ;
        RECT 343.810 395.720 365.050 396.000 ;
        RECT 365.890 395.720 387.130 396.000 ;
        RECT 12.060 10.695 387.680 395.720 ;
      LAYER met3 ;
        RECT 21.050 10.715 329.830 389.125 ;
  END
END arbiterpuf
END LIBRARY

