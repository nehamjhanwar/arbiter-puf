magic
tech sky130A
magscale 1 2
timestamp 1671600370
<< nwell >>
rect 1066 77509 78882 77830
rect 1066 76421 78882 76987
rect 1066 75333 78882 75899
rect 1066 74245 78882 74811
rect 1066 73157 78882 73723
rect 1066 72069 78882 72635
rect 1066 70981 78882 71547
rect 1066 69893 78882 70459
rect 1066 68805 78882 69371
rect 1066 67717 78882 68283
rect 1066 66629 78882 67195
rect 1066 65541 78882 66107
rect 1066 64453 78882 65019
rect 1066 63365 78882 63931
rect 1066 62277 78882 62843
rect 1066 61189 78882 61755
rect 1066 60101 78882 60667
rect 1066 59013 78882 59579
rect 1066 57925 78882 58491
rect 1066 56837 78882 57403
rect 1066 55749 78882 56315
rect 1066 54661 78882 55227
rect 1066 53573 78882 54139
rect 1066 52485 78882 53051
rect 1066 51397 78882 51963
rect 1066 50309 78882 50875
rect 1066 49221 78882 49787
rect 1066 48133 78882 48699
rect 1066 47045 78882 47611
rect 1066 45957 78882 46523
rect 1066 44869 78882 45435
rect 1066 43781 78882 44347
rect 1066 42693 78882 43259
rect 1066 41605 78882 42171
rect 1066 40517 78882 41083
rect 1066 39429 78882 39995
rect 1066 38341 78882 38907
rect 1066 37253 78882 37819
rect 1066 36165 78882 36731
rect 1066 35077 78882 35643
rect 1066 33989 78882 34555
rect 1066 32901 78882 33467
rect 1066 31813 78882 32379
rect 1066 30725 78882 31291
rect 1066 29637 78882 30203
rect 1066 28549 78882 29115
rect 1066 27461 78882 28027
rect 1066 26373 78882 26939
rect 1066 25285 78882 25851
rect 1066 24197 78882 24763
rect 1066 23109 78882 23675
rect 1066 22021 78882 22587
rect 1066 20933 78882 21499
rect 1066 19845 78882 20411
rect 1066 18757 78882 19323
rect 1066 17669 78882 18235
rect 1066 16581 78882 17147
rect 1066 15493 78882 16059
rect 1066 14405 78882 14971
rect 1066 13317 78882 13883
rect 1066 12229 78882 12795
rect 1066 11141 78882 11707
rect 1066 10053 78882 10619
rect 1066 8965 78882 9531
rect 1066 7877 78882 8443
rect 1066 6789 78882 7355
rect 1066 5701 78882 6267
rect 1066 4613 78882 5179
rect 1066 3525 78882 4091
rect 1066 2437 78882 3003
<< obsli1 >>
rect 1104 2159 78844 77809
<< obsm1 >>
rect 1104 2128 78844 77840
<< metal2 >>
rect 2410 79200 2466 80000
rect 6826 79200 6882 80000
rect 11242 79200 11298 80000
rect 15658 79200 15714 80000
rect 20074 79200 20130 80000
rect 24490 79200 24546 80000
rect 28906 79200 28962 80000
rect 33322 79200 33378 80000
rect 37738 79200 37794 80000
rect 42154 79200 42210 80000
rect 46570 79200 46626 80000
rect 50986 79200 51042 80000
rect 55402 79200 55458 80000
rect 59818 79200 59874 80000
rect 64234 79200 64290 80000
rect 68650 79200 68706 80000
rect 73066 79200 73122 80000
rect 77482 79200 77538 80000
<< obsm2 >>
rect 2522 79144 6770 79200
rect 6938 79144 11186 79200
rect 11354 79144 15602 79200
rect 15770 79144 20018 79200
rect 20186 79144 24434 79200
rect 24602 79144 28850 79200
rect 29018 79144 33266 79200
rect 33434 79144 37682 79200
rect 37850 79144 42098 79200
rect 42266 79144 46514 79200
rect 46682 79144 50930 79200
rect 51098 79144 55346 79200
rect 55514 79144 59762 79200
rect 59930 79144 64178 79200
rect 64346 79144 68594 79200
rect 68762 79144 73010 79200
rect 73178 79144 77426 79200
rect 2412 2139 77536 79144
<< obsm3 >>
rect 4210 2143 65966 77825
<< metal4 >>
rect 4208 2128 4528 77840
rect 19568 2128 19888 77840
rect 34928 2128 35248 77840
rect 50288 2128 50608 77840
rect 65648 2128 65968 77840
<< labels >>
rlabel metal2 s 6826 79200 6882 80000 6 ichallenge[0]
port 1 nsew signal input
rlabel metal2 s 50986 79200 51042 80000 6 ichallenge[10]
port 2 nsew signal input
rlabel metal2 s 55402 79200 55458 80000 6 ichallenge[11]
port 3 nsew signal input
rlabel metal2 s 59818 79200 59874 80000 6 ichallenge[12]
port 4 nsew signal input
rlabel metal2 s 64234 79200 64290 80000 6 ichallenge[13]
port 5 nsew signal input
rlabel metal2 s 68650 79200 68706 80000 6 ichallenge[14]
port 6 nsew signal input
rlabel metal2 s 73066 79200 73122 80000 6 ichallenge[15]
port 7 nsew signal input
rlabel metal2 s 11242 79200 11298 80000 6 ichallenge[1]
port 8 nsew signal input
rlabel metal2 s 15658 79200 15714 80000 6 ichallenge[2]
port 9 nsew signal input
rlabel metal2 s 20074 79200 20130 80000 6 ichallenge[3]
port 10 nsew signal input
rlabel metal2 s 24490 79200 24546 80000 6 ichallenge[4]
port 11 nsew signal input
rlabel metal2 s 28906 79200 28962 80000 6 ichallenge[5]
port 12 nsew signal input
rlabel metal2 s 33322 79200 33378 80000 6 ichallenge[6]
port 13 nsew signal input
rlabel metal2 s 37738 79200 37794 80000 6 ichallenge[7]
port 14 nsew signal input
rlabel metal2 s 42154 79200 42210 80000 6 ichallenge[8]
port 15 nsew signal input
rlabel metal2 s 46570 79200 46626 80000 6 ichallenge[9]
port 16 nsew signal input
rlabel metal2 s 2410 79200 2466 80000 6 ipulse
port 17 nsew signal input
rlabel metal2 s 77482 79200 77538 80000 6 oresponse
port 18 nsew signal output
rlabel metal4 s 4208 2128 4528 77840 6 vccd1
port 19 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 77840 6 vccd1
port 19 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 77840 6 vccd1
port 19 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 77840 6 vssd1
port 20 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 77840 6 vssd1
port 20 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 80000 80000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 1587926
string GDS_FILE /home/radhe/project/matrix_multiply_mpw8/openlane/arbiterpuf/runs/22_12_21_10_47/results/signoff/arbiterpuf.magic.gds
string GDS_START 45102
<< end >>

