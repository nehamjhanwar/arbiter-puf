magic
tech sky130A
magscale 1 2
timestamp 1671452076
<< nwell >>
rect 1066 116677 178886 117243
rect 1066 115589 178886 116155
rect 1066 114501 178886 115067
rect 1066 113413 178886 113979
rect 1066 112325 178886 112891
rect 1066 111237 178886 111803
rect 1066 110149 178886 110715
rect 1066 109061 178886 109627
rect 1066 107973 178886 108539
rect 1066 106885 178886 107451
rect 1066 105797 178886 106363
rect 1066 104709 178886 105275
rect 1066 103621 178886 104187
rect 1066 102533 178886 103099
rect 1066 101445 178886 102011
rect 1066 100357 178886 100923
rect 1066 99269 178886 99835
rect 1066 98181 178886 98747
rect 1066 97093 178886 97659
rect 1066 96005 178886 96571
rect 1066 94917 178886 95483
rect 1066 93829 178886 94395
rect 1066 92741 178886 93307
rect 1066 91653 178886 92219
rect 1066 90565 178886 91131
rect 1066 89477 178886 90043
rect 1066 88389 178886 88955
rect 1066 87301 178886 87867
rect 1066 86213 178886 86779
rect 1066 85125 178886 85691
rect 1066 84037 178886 84603
rect 1066 82949 178886 83515
rect 1066 81861 178886 82427
rect 1066 80773 178886 81339
rect 1066 79685 178886 80251
rect 1066 78597 178886 79163
rect 1066 77509 178886 78075
rect 1066 76421 178886 76987
rect 1066 75333 178886 75899
rect 1066 74245 178886 74811
rect 1066 73157 178886 73723
rect 1066 72069 178886 72635
rect 1066 70981 178886 71547
rect 1066 69893 178886 70459
rect 1066 68805 178886 69371
rect 1066 67717 178886 68283
rect 1066 66629 178886 67195
rect 1066 65541 178886 66107
rect 1066 64453 178886 65019
rect 1066 63365 178886 63931
rect 1066 62277 178886 62843
rect 1066 61189 178886 61755
rect 1066 60101 178886 60667
rect 1066 59013 178886 59579
rect 1066 57925 178886 58491
rect 1066 56837 178886 57403
rect 1066 55749 178886 56315
rect 1066 54661 178886 55227
rect 1066 53573 178886 54139
rect 1066 52485 178886 53051
rect 1066 51397 178886 51963
rect 1066 50309 178886 50875
rect 1066 49221 178886 49787
rect 1066 48133 178886 48699
rect 1066 47045 178886 47611
rect 1066 45957 178886 46523
rect 1066 44869 178886 45435
rect 1066 43781 178886 44347
rect 1066 42693 178886 43259
rect 1066 41605 178886 42171
rect 1066 40517 178886 41083
rect 1066 39429 178886 39995
rect 1066 38341 178886 38907
rect 1066 37253 178886 37819
rect 1066 36165 178886 36731
rect 1066 35077 178886 35643
rect 1066 33989 178886 34555
rect 1066 32901 178886 33467
rect 1066 31813 178886 32379
rect 1066 30725 178886 31291
rect 1066 29637 178886 30203
rect 1066 28549 178886 29115
rect 1066 27461 178886 28027
rect 1066 26373 178886 26939
rect 1066 25285 178886 25851
rect 1066 24197 178886 24763
rect 1066 23109 178886 23675
rect 1066 22021 178886 22587
rect 1066 20933 178886 21499
rect 1066 19845 178886 20411
rect 1066 18757 178886 19323
rect 1066 17669 178886 18235
rect 1066 16581 178886 17147
rect 1066 15493 178886 16059
rect 1066 14405 178886 14971
rect 1066 13317 178886 13883
rect 1066 12229 178886 12795
rect 1066 11141 178886 11707
rect 1066 10053 178886 10619
rect 1066 8965 178886 9531
rect 1066 7877 178886 8443
rect 1066 6789 178886 7355
rect 1066 5701 178886 6267
rect 1066 4613 178886 5179
rect 1066 3525 178886 4091
rect 1066 2437 178886 3003
<< obsli1 >>
rect 1104 2159 178848 117521
<< obsm1 >>
rect 1104 1436 178848 117552
<< metal2 >>
rect 3054 0 3110 800
rect 8482 0 8538 800
rect 13910 0 13966 800
rect 19338 0 19394 800
rect 24766 0 24822 800
rect 30194 0 30250 800
rect 35622 0 35678 800
rect 41050 0 41106 800
rect 46478 0 46534 800
rect 51906 0 51962 800
rect 57334 0 57390 800
rect 62762 0 62818 800
rect 68190 0 68246 800
rect 73618 0 73674 800
rect 79046 0 79102 800
rect 84474 0 84530 800
rect 89902 0 89958 800
rect 95330 0 95386 800
rect 100758 0 100814 800
rect 106186 0 106242 800
rect 111614 0 111670 800
rect 117042 0 117098 800
rect 122470 0 122526 800
rect 127898 0 127954 800
rect 133326 0 133382 800
rect 138754 0 138810 800
rect 144182 0 144238 800
rect 149610 0 149666 800
rect 155038 0 155094 800
rect 160466 0 160522 800
rect 165894 0 165950 800
rect 171322 0 171378 800
rect 176750 0 176806 800
<< obsm2 >>
rect 3056 856 176804 117541
rect 3166 800 8426 856
rect 8594 800 13854 856
rect 14022 800 19282 856
rect 19450 800 24710 856
rect 24878 800 30138 856
rect 30306 800 35566 856
rect 35734 800 40994 856
rect 41162 800 46422 856
rect 46590 800 51850 856
rect 52018 800 57278 856
rect 57446 800 62706 856
rect 62874 800 68134 856
rect 68302 800 73562 856
rect 73730 800 78990 856
rect 79158 800 84418 856
rect 84586 800 89846 856
rect 90014 800 95274 856
rect 95442 800 100702 856
rect 100870 800 106130 856
rect 106298 800 111558 856
rect 111726 800 116986 856
rect 117154 800 122414 856
rect 122582 800 127842 856
rect 128010 800 133270 856
rect 133438 800 138698 856
rect 138866 800 144126 856
rect 144294 800 149554 856
rect 149722 800 154982 856
rect 155150 800 160410 856
rect 160578 800 165838 856
rect 166006 800 171266 856
rect 171434 800 176694 856
<< obsm3 >>
rect 4153 2143 176719 117537
<< metal4 >>
rect 4208 2128 4528 117552
rect 19568 2128 19888 117552
rect 34928 2128 35248 117552
rect 50288 2128 50608 117552
rect 65648 2128 65968 117552
rect 81008 2128 81328 117552
rect 96368 2128 96688 117552
rect 111728 2128 112048 117552
rect 127088 2128 127408 117552
rect 142448 2128 142768 117552
rect 157808 2128 158128 117552
rect 173168 2128 173488 117552
<< obsm4 >>
rect 11651 2211 19488 34917
rect 19968 2211 34848 34917
rect 35328 2211 50208 34917
rect 50688 2211 65568 34917
rect 66048 2211 80928 34917
rect 81408 2211 88445 34917
<< labels >>
rlabel metal2 s 13910 0 13966 800 6 clk
port 1 nsew signal input
rlabel metal2 s 8482 0 8538 800 6 execute
port 2 nsew signal input
rlabel metal2 s 35622 0 35678 800 6 input_val[0]
port 3 nsew signal input
rlabel metal2 s 41050 0 41106 800 6 input_val[1]
port 4 nsew signal input
rlabel metal2 s 46478 0 46534 800 6 input_val[2]
port 5 nsew signal input
rlabel metal2 s 51906 0 51962 800 6 input_val[3]
port 6 nsew signal input
rlabel metal2 s 57334 0 57390 800 6 input_val[4]
port 7 nsew signal input
rlabel metal2 s 62762 0 62818 800 6 input_val[5]
port 8 nsew signal input
rlabel metal2 s 68190 0 68246 800 6 input_val[6]
port 9 nsew signal input
rlabel metal2 s 73618 0 73674 800 6 input_val[7]
port 10 nsew signal input
rlabel metal2 s 3054 0 3110 800 6 reset
port 11 nsew signal input
rlabel metal2 s 89902 0 89958 800 6 result[0]
port 12 nsew signal output
rlabel metal2 s 144182 0 144238 800 6 result[10]
port 13 nsew signal output
rlabel metal2 s 149610 0 149666 800 6 result[11]
port 14 nsew signal output
rlabel metal2 s 155038 0 155094 800 6 result[12]
port 15 nsew signal output
rlabel metal2 s 160466 0 160522 800 6 result[13]
port 16 nsew signal output
rlabel metal2 s 165894 0 165950 800 6 result[14]
port 17 nsew signal output
rlabel metal2 s 171322 0 171378 800 6 result[15]
port 18 nsew signal output
rlabel metal2 s 176750 0 176806 800 6 result[16]
port 19 nsew signal output
rlabel metal2 s 95330 0 95386 800 6 result[1]
port 20 nsew signal output
rlabel metal2 s 100758 0 100814 800 6 result[2]
port 21 nsew signal output
rlabel metal2 s 106186 0 106242 800 6 result[3]
port 22 nsew signal output
rlabel metal2 s 111614 0 111670 800 6 result[4]
port 23 nsew signal output
rlabel metal2 s 117042 0 117098 800 6 result[5]
port 24 nsew signal output
rlabel metal2 s 122470 0 122526 800 6 result[6]
port 25 nsew signal output
rlabel metal2 s 127898 0 127954 800 6 result[7]
port 26 nsew signal output
rlabel metal2 s 133326 0 133382 800 6 result[8]
port 27 nsew signal output
rlabel metal2 s 138754 0 138810 800 6 result[9]
port 28 nsew signal output
rlabel metal2 s 19338 0 19394 800 6 sel_in[0]
port 29 nsew signal input
rlabel metal2 s 24766 0 24822 800 6 sel_in[1]
port 30 nsew signal input
rlabel metal2 s 30194 0 30250 800 6 sel_in[2]
port 31 nsew signal input
rlabel metal2 s 79046 0 79102 800 6 sel_out[0]
port 32 nsew signal input
rlabel metal2 s 84474 0 84530 800 6 sel_out[1]
port 33 nsew signal input
rlabel metal4 s 4208 2128 4528 117552 6 vccd1
port 34 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 117552 6 vccd1
port 34 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 117552 6 vccd1
port 34 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 117552 6 vccd1
port 34 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 117552 6 vccd1
port 34 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 117552 6 vccd1
port 34 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 117552 6 vssd1
port 35 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 117552 6 vssd1
port 35 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 117552 6 vssd1
port 35 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 117552 6 vssd1
port 35 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 117552 6 vssd1
port 35 nsew ground bidirectional
rlabel metal4 s 173168 2128 173488 117552 6 vssd1
port 35 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 180000 120000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 16243594
string GDS_FILE /home/radhe/project/matrix_multiply_mpw8/openlane/matrix_multiply/runs/22_12_19_16_52/results/signoff/matrix_multiply.magic.gds
string GDS_START 845128
<< end >>

