magic
tech sky130A
magscale 1 2
timestamp 1671356593
<< obsli1 >>
rect 1104 2159 178848 117521
<< obsm1 >>
rect 1104 2128 178848 117552
<< metal2 >>
rect 3790 119200 3846 120000
rect 10414 119200 10470 120000
rect 17038 119200 17094 120000
rect 23662 119200 23718 120000
rect 30286 119200 30342 120000
rect 36910 119200 36966 120000
rect 43534 119200 43590 120000
rect 50158 119200 50214 120000
rect 56782 119200 56838 120000
rect 63406 119200 63462 120000
rect 70030 119200 70086 120000
rect 76654 119200 76710 120000
rect 83278 119200 83334 120000
rect 89902 119200 89958 120000
rect 96526 119200 96582 120000
rect 103150 119200 103206 120000
rect 109774 119200 109830 120000
rect 116398 119200 116454 120000
rect 123022 119200 123078 120000
rect 129646 119200 129702 120000
rect 136270 119200 136326 120000
rect 142894 119200 142950 120000
rect 149518 119200 149574 120000
rect 156142 119200 156198 120000
rect 162766 119200 162822 120000
rect 169390 119200 169446 120000
rect 176014 119200 176070 120000
rect 6826 0 6882 800
rect 7378 0 7434 800
rect 7930 0 7986 800
rect 8482 0 8538 800
rect 9034 0 9090 800
rect 9586 0 9642 800
rect 10138 0 10194 800
rect 10690 0 10746 800
rect 11242 0 11298 800
rect 11794 0 11850 800
rect 12346 0 12402 800
rect 12898 0 12954 800
rect 13450 0 13506 800
rect 14002 0 14058 800
rect 14554 0 14610 800
rect 15106 0 15162 800
rect 15658 0 15714 800
rect 16210 0 16266 800
rect 16762 0 16818 800
rect 17314 0 17370 800
rect 17866 0 17922 800
rect 18418 0 18474 800
rect 18970 0 19026 800
rect 19522 0 19578 800
rect 20074 0 20130 800
rect 20626 0 20682 800
rect 21178 0 21234 800
rect 21730 0 21786 800
rect 22282 0 22338 800
rect 22834 0 22890 800
rect 23386 0 23442 800
rect 23938 0 23994 800
rect 24490 0 24546 800
rect 25042 0 25098 800
rect 25594 0 25650 800
rect 26146 0 26202 800
rect 26698 0 26754 800
rect 27250 0 27306 800
rect 27802 0 27858 800
rect 28354 0 28410 800
rect 28906 0 28962 800
rect 29458 0 29514 800
rect 30010 0 30066 800
rect 30562 0 30618 800
rect 31114 0 31170 800
rect 31666 0 31722 800
rect 32218 0 32274 800
rect 32770 0 32826 800
rect 33322 0 33378 800
rect 33874 0 33930 800
rect 34426 0 34482 800
rect 34978 0 35034 800
rect 35530 0 35586 800
rect 36082 0 36138 800
rect 36634 0 36690 800
rect 37186 0 37242 800
rect 37738 0 37794 800
rect 38290 0 38346 800
rect 38842 0 38898 800
rect 39394 0 39450 800
rect 39946 0 40002 800
rect 40498 0 40554 800
rect 41050 0 41106 800
rect 41602 0 41658 800
rect 42154 0 42210 800
rect 42706 0 42762 800
rect 43258 0 43314 800
rect 43810 0 43866 800
rect 44362 0 44418 800
rect 44914 0 44970 800
rect 45466 0 45522 800
rect 46018 0 46074 800
rect 46570 0 46626 800
rect 47122 0 47178 800
rect 47674 0 47730 800
rect 48226 0 48282 800
rect 48778 0 48834 800
rect 49330 0 49386 800
rect 49882 0 49938 800
rect 50434 0 50490 800
rect 50986 0 51042 800
rect 51538 0 51594 800
rect 52090 0 52146 800
rect 52642 0 52698 800
rect 53194 0 53250 800
rect 53746 0 53802 800
rect 54298 0 54354 800
rect 54850 0 54906 800
rect 55402 0 55458 800
rect 55954 0 56010 800
rect 56506 0 56562 800
rect 57058 0 57114 800
rect 57610 0 57666 800
rect 58162 0 58218 800
rect 58714 0 58770 800
rect 59266 0 59322 800
rect 59818 0 59874 800
rect 60370 0 60426 800
rect 60922 0 60978 800
rect 61474 0 61530 800
rect 62026 0 62082 800
rect 62578 0 62634 800
rect 63130 0 63186 800
rect 63682 0 63738 800
rect 64234 0 64290 800
rect 64786 0 64842 800
rect 65338 0 65394 800
rect 65890 0 65946 800
rect 66442 0 66498 800
rect 66994 0 67050 800
rect 67546 0 67602 800
rect 68098 0 68154 800
rect 68650 0 68706 800
rect 69202 0 69258 800
rect 69754 0 69810 800
rect 70306 0 70362 800
rect 70858 0 70914 800
rect 71410 0 71466 800
rect 71962 0 72018 800
rect 72514 0 72570 800
rect 73066 0 73122 800
rect 73618 0 73674 800
rect 74170 0 74226 800
rect 74722 0 74778 800
rect 75274 0 75330 800
rect 75826 0 75882 800
rect 76378 0 76434 800
rect 76930 0 76986 800
rect 77482 0 77538 800
rect 78034 0 78090 800
rect 78586 0 78642 800
rect 79138 0 79194 800
rect 79690 0 79746 800
rect 80242 0 80298 800
rect 80794 0 80850 800
rect 81346 0 81402 800
rect 81898 0 81954 800
rect 82450 0 82506 800
rect 83002 0 83058 800
rect 83554 0 83610 800
rect 84106 0 84162 800
rect 84658 0 84714 800
rect 85210 0 85266 800
rect 85762 0 85818 800
rect 86314 0 86370 800
rect 86866 0 86922 800
rect 87418 0 87474 800
rect 87970 0 88026 800
rect 88522 0 88578 800
rect 89074 0 89130 800
rect 89626 0 89682 800
rect 90178 0 90234 800
rect 90730 0 90786 800
rect 91282 0 91338 800
rect 91834 0 91890 800
rect 92386 0 92442 800
rect 92938 0 92994 800
rect 93490 0 93546 800
rect 94042 0 94098 800
rect 94594 0 94650 800
rect 95146 0 95202 800
rect 95698 0 95754 800
rect 96250 0 96306 800
rect 96802 0 96858 800
rect 97354 0 97410 800
rect 97906 0 97962 800
rect 98458 0 98514 800
rect 99010 0 99066 800
rect 99562 0 99618 800
rect 100114 0 100170 800
rect 100666 0 100722 800
rect 101218 0 101274 800
rect 101770 0 101826 800
rect 102322 0 102378 800
rect 102874 0 102930 800
rect 103426 0 103482 800
rect 103978 0 104034 800
rect 104530 0 104586 800
rect 105082 0 105138 800
rect 105634 0 105690 800
rect 106186 0 106242 800
rect 106738 0 106794 800
rect 107290 0 107346 800
rect 107842 0 107898 800
rect 108394 0 108450 800
rect 108946 0 109002 800
rect 109498 0 109554 800
rect 110050 0 110106 800
rect 110602 0 110658 800
rect 111154 0 111210 800
rect 111706 0 111762 800
rect 112258 0 112314 800
rect 112810 0 112866 800
rect 113362 0 113418 800
rect 113914 0 113970 800
rect 114466 0 114522 800
rect 115018 0 115074 800
rect 115570 0 115626 800
rect 116122 0 116178 800
rect 116674 0 116730 800
rect 117226 0 117282 800
rect 117778 0 117834 800
rect 118330 0 118386 800
rect 118882 0 118938 800
rect 119434 0 119490 800
rect 119986 0 120042 800
rect 120538 0 120594 800
rect 121090 0 121146 800
rect 121642 0 121698 800
rect 122194 0 122250 800
rect 122746 0 122802 800
rect 123298 0 123354 800
rect 123850 0 123906 800
rect 124402 0 124458 800
rect 124954 0 125010 800
rect 125506 0 125562 800
rect 126058 0 126114 800
rect 126610 0 126666 800
rect 127162 0 127218 800
rect 127714 0 127770 800
rect 128266 0 128322 800
rect 128818 0 128874 800
rect 129370 0 129426 800
rect 129922 0 129978 800
rect 130474 0 130530 800
rect 131026 0 131082 800
rect 131578 0 131634 800
rect 132130 0 132186 800
rect 132682 0 132738 800
rect 133234 0 133290 800
rect 133786 0 133842 800
rect 134338 0 134394 800
rect 134890 0 134946 800
rect 135442 0 135498 800
rect 135994 0 136050 800
rect 136546 0 136602 800
rect 137098 0 137154 800
rect 137650 0 137706 800
rect 138202 0 138258 800
rect 138754 0 138810 800
rect 139306 0 139362 800
rect 139858 0 139914 800
rect 140410 0 140466 800
rect 140962 0 141018 800
rect 141514 0 141570 800
rect 142066 0 142122 800
rect 142618 0 142674 800
rect 143170 0 143226 800
rect 143722 0 143778 800
rect 144274 0 144330 800
rect 144826 0 144882 800
rect 145378 0 145434 800
rect 145930 0 145986 800
rect 146482 0 146538 800
rect 147034 0 147090 800
rect 147586 0 147642 800
rect 148138 0 148194 800
rect 148690 0 148746 800
rect 149242 0 149298 800
rect 149794 0 149850 800
rect 150346 0 150402 800
rect 150898 0 150954 800
rect 151450 0 151506 800
rect 152002 0 152058 800
rect 152554 0 152610 800
rect 153106 0 153162 800
rect 153658 0 153714 800
rect 154210 0 154266 800
rect 154762 0 154818 800
rect 155314 0 155370 800
rect 155866 0 155922 800
rect 156418 0 156474 800
rect 156970 0 157026 800
rect 157522 0 157578 800
rect 158074 0 158130 800
rect 158626 0 158682 800
rect 159178 0 159234 800
rect 159730 0 159786 800
rect 160282 0 160338 800
rect 160834 0 160890 800
rect 161386 0 161442 800
rect 161938 0 161994 800
rect 162490 0 162546 800
rect 163042 0 163098 800
rect 163594 0 163650 800
rect 164146 0 164202 800
rect 164698 0 164754 800
rect 165250 0 165306 800
rect 165802 0 165858 800
rect 166354 0 166410 800
rect 166906 0 166962 800
rect 167458 0 167514 800
rect 168010 0 168066 800
rect 168562 0 168618 800
rect 169114 0 169170 800
rect 169666 0 169722 800
rect 170218 0 170274 800
rect 170770 0 170826 800
rect 171322 0 171378 800
rect 171874 0 171930 800
rect 172426 0 172482 800
rect 172978 0 173034 800
<< obsm2 >>
rect 1582 119144 3734 119354
rect 3902 119144 10358 119354
rect 10526 119144 16982 119354
rect 17150 119144 23606 119354
rect 23774 119144 30230 119354
rect 30398 119144 36854 119354
rect 37022 119144 43478 119354
rect 43646 119144 50102 119354
rect 50270 119144 56726 119354
rect 56894 119144 63350 119354
rect 63518 119144 69974 119354
rect 70142 119144 76598 119354
rect 76766 119144 83222 119354
rect 83390 119144 89846 119354
rect 90014 119144 96470 119354
rect 96638 119144 103094 119354
rect 103262 119144 109718 119354
rect 109886 119144 116342 119354
rect 116510 119144 122966 119354
rect 123134 119144 129590 119354
rect 129758 119144 136214 119354
rect 136382 119144 142838 119354
rect 143006 119144 149462 119354
rect 149630 119144 156086 119354
rect 156254 119144 162710 119354
rect 162878 119144 169334 119354
rect 169502 119144 175958 119354
rect 176126 119144 178370 119354
rect 1582 856 178370 119144
rect 1582 800 6770 856
rect 6938 800 7322 856
rect 7490 800 7874 856
rect 8042 800 8426 856
rect 8594 800 8978 856
rect 9146 800 9530 856
rect 9698 800 10082 856
rect 10250 800 10634 856
rect 10802 800 11186 856
rect 11354 800 11738 856
rect 11906 800 12290 856
rect 12458 800 12842 856
rect 13010 800 13394 856
rect 13562 800 13946 856
rect 14114 800 14498 856
rect 14666 800 15050 856
rect 15218 800 15602 856
rect 15770 800 16154 856
rect 16322 800 16706 856
rect 16874 800 17258 856
rect 17426 800 17810 856
rect 17978 800 18362 856
rect 18530 800 18914 856
rect 19082 800 19466 856
rect 19634 800 20018 856
rect 20186 800 20570 856
rect 20738 800 21122 856
rect 21290 800 21674 856
rect 21842 800 22226 856
rect 22394 800 22778 856
rect 22946 800 23330 856
rect 23498 800 23882 856
rect 24050 800 24434 856
rect 24602 800 24986 856
rect 25154 800 25538 856
rect 25706 800 26090 856
rect 26258 800 26642 856
rect 26810 800 27194 856
rect 27362 800 27746 856
rect 27914 800 28298 856
rect 28466 800 28850 856
rect 29018 800 29402 856
rect 29570 800 29954 856
rect 30122 800 30506 856
rect 30674 800 31058 856
rect 31226 800 31610 856
rect 31778 800 32162 856
rect 32330 800 32714 856
rect 32882 800 33266 856
rect 33434 800 33818 856
rect 33986 800 34370 856
rect 34538 800 34922 856
rect 35090 800 35474 856
rect 35642 800 36026 856
rect 36194 800 36578 856
rect 36746 800 37130 856
rect 37298 800 37682 856
rect 37850 800 38234 856
rect 38402 800 38786 856
rect 38954 800 39338 856
rect 39506 800 39890 856
rect 40058 800 40442 856
rect 40610 800 40994 856
rect 41162 800 41546 856
rect 41714 800 42098 856
rect 42266 800 42650 856
rect 42818 800 43202 856
rect 43370 800 43754 856
rect 43922 800 44306 856
rect 44474 800 44858 856
rect 45026 800 45410 856
rect 45578 800 45962 856
rect 46130 800 46514 856
rect 46682 800 47066 856
rect 47234 800 47618 856
rect 47786 800 48170 856
rect 48338 800 48722 856
rect 48890 800 49274 856
rect 49442 800 49826 856
rect 49994 800 50378 856
rect 50546 800 50930 856
rect 51098 800 51482 856
rect 51650 800 52034 856
rect 52202 800 52586 856
rect 52754 800 53138 856
rect 53306 800 53690 856
rect 53858 800 54242 856
rect 54410 800 54794 856
rect 54962 800 55346 856
rect 55514 800 55898 856
rect 56066 800 56450 856
rect 56618 800 57002 856
rect 57170 800 57554 856
rect 57722 800 58106 856
rect 58274 800 58658 856
rect 58826 800 59210 856
rect 59378 800 59762 856
rect 59930 800 60314 856
rect 60482 800 60866 856
rect 61034 800 61418 856
rect 61586 800 61970 856
rect 62138 800 62522 856
rect 62690 800 63074 856
rect 63242 800 63626 856
rect 63794 800 64178 856
rect 64346 800 64730 856
rect 64898 800 65282 856
rect 65450 800 65834 856
rect 66002 800 66386 856
rect 66554 800 66938 856
rect 67106 800 67490 856
rect 67658 800 68042 856
rect 68210 800 68594 856
rect 68762 800 69146 856
rect 69314 800 69698 856
rect 69866 800 70250 856
rect 70418 800 70802 856
rect 70970 800 71354 856
rect 71522 800 71906 856
rect 72074 800 72458 856
rect 72626 800 73010 856
rect 73178 800 73562 856
rect 73730 800 74114 856
rect 74282 800 74666 856
rect 74834 800 75218 856
rect 75386 800 75770 856
rect 75938 800 76322 856
rect 76490 800 76874 856
rect 77042 800 77426 856
rect 77594 800 77978 856
rect 78146 800 78530 856
rect 78698 800 79082 856
rect 79250 800 79634 856
rect 79802 800 80186 856
rect 80354 800 80738 856
rect 80906 800 81290 856
rect 81458 800 81842 856
rect 82010 800 82394 856
rect 82562 800 82946 856
rect 83114 800 83498 856
rect 83666 800 84050 856
rect 84218 800 84602 856
rect 84770 800 85154 856
rect 85322 800 85706 856
rect 85874 800 86258 856
rect 86426 800 86810 856
rect 86978 800 87362 856
rect 87530 800 87914 856
rect 88082 800 88466 856
rect 88634 800 89018 856
rect 89186 800 89570 856
rect 89738 800 90122 856
rect 90290 800 90674 856
rect 90842 800 91226 856
rect 91394 800 91778 856
rect 91946 800 92330 856
rect 92498 800 92882 856
rect 93050 800 93434 856
rect 93602 800 93986 856
rect 94154 800 94538 856
rect 94706 800 95090 856
rect 95258 800 95642 856
rect 95810 800 96194 856
rect 96362 800 96746 856
rect 96914 800 97298 856
rect 97466 800 97850 856
rect 98018 800 98402 856
rect 98570 800 98954 856
rect 99122 800 99506 856
rect 99674 800 100058 856
rect 100226 800 100610 856
rect 100778 800 101162 856
rect 101330 800 101714 856
rect 101882 800 102266 856
rect 102434 800 102818 856
rect 102986 800 103370 856
rect 103538 800 103922 856
rect 104090 800 104474 856
rect 104642 800 105026 856
rect 105194 800 105578 856
rect 105746 800 106130 856
rect 106298 800 106682 856
rect 106850 800 107234 856
rect 107402 800 107786 856
rect 107954 800 108338 856
rect 108506 800 108890 856
rect 109058 800 109442 856
rect 109610 800 109994 856
rect 110162 800 110546 856
rect 110714 800 111098 856
rect 111266 800 111650 856
rect 111818 800 112202 856
rect 112370 800 112754 856
rect 112922 800 113306 856
rect 113474 800 113858 856
rect 114026 800 114410 856
rect 114578 800 114962 856
rect 115130 800 115514 856
rect 115682 800 116066 856
rect 116234 800 116618 856
rect 116786 800 117170 856
rect 117338 800 117722 856
rect 117890 800 118274 856
rect 118442 800 118826 856
rect 118994 800 119378 856
rect 119546 800 119930 856
rect 120098 800 120482 856
rect 120650 800 121034 856
rect 121202 800 121586 856
rect 121754 800 122138 856
rect 122306 800 122690 856
rect 122858 800 123242 856
rect 123410 800 123794 856
rect 123962 800 124346 856
rect 124514 800 124898 856
rect 125066 800 125450 856
rect 125618 800 126002 856
rect 126170 800 126554 856
rect 126722 800 127106 856
rect 127274 800 127658 856
rect 127826 800 128210 856
rect 128378 800 128762 856
rect 128930 800 129314 856
rect 129482 800 129866 856
rect 130034 800 130418 856
rect 130586 800 130970 856
rect 131138 800 131522 856
rect 131690 800 132074 856
rect 132242 800 132626 856
rect 132794 800 133178 856
rect 133346 800 133730 856
rect 133898 800 134282 856
rect 134450 800 134834 856
rect 135002 800 135386 856
rect 135554 800 135938 856
rect 136106 800 136490 856
rect 136658 800 137042 856
rect 137210 800 137594 856
rect 137762 800 138146 856
rect 138314 800 138698 856
rect 138866 800 139250 856
rect 139418 800 139802 856
rect 139970 800 140354 856
rect 140522 800 140906 856
rect 141074 800 141458 856
rect 141626 800 142010 856
rect 142178 800 142562 856
rect 142730 800 143114 856
rect 143282 800 143666 856
rect 143834 800 144218 856
rect 144386 800 144770 856
rect 144938 800 145322 856
rect 145490 800 145874 856
rect 146042 800 146426 856
rect 146594 800 146978 856
rect 147146 800 147530 856
rect 147698 800 148082 856
rect 148250 800 148634 856
rect 148802 800 149186 856
rect 149354 800 149738 856
rect 149906 800 150290 856
rect 150458 800 150842 856
rect 151010 800 151394 856
rect 151562 800 151946 856
rect 152114 800 152498 856
rect 152666 800 153050 856
rect 153218 800 153602 856
rect 153770 800 154154 856
rect 154322 800 154706 856
rect 154874 800 155258 856
rect 155426 800 155810 856
rect 155978 800 156362 856
rect 156530 800 156914 856
rect 157082 800 157466 856
rect 157634 800 158018 856
rect 158186 800 158570 856
rect 158738 800 159122 856
rect 159290 800 159674 856
rect 159842 800 160226 856
rect 160394 800 160778 856
rect 160946 800 161330 856
rect 161498 800 161882 856
rect 162050 800 162434 856
rect 162602 800 162986 856
rect 163154 800 163538 856
rect 163706 800 164090 856
rect 164258 800 164642 856
rect 164810 800 165194 856
rect 165362 800 165746 856
rect 165914 800 166298 856
rect 166466 800 166850 856
rect 167018 800 167402 856
rect 167570 800 167954 856
rect 168122 800 168506 856
rect 168674 800 169058 856
rect 169226 800 169610 856
rect 169778 800 170162 856
rect 170330 800 170714 856
rect 170882 800 171266 856
rect 171434 800 171818 856
rect 171986 800 172370 856
rect 172538 800 172922 856
rect 173090 800 178370 856
<< metal3 >>
rect 0 118464 800 118584
rect 179200 116696 180000 116816
rect 0 115608 800 115728
rect 179200 114112 180000 114232
rect 0 112752 800 112872
rect 179200 111528 180000 111648
rect 0 109896 800 110016
rect 179200 108944 180000 109064
rect 0 107040 800 107160
rect 179200 106360 180000 106480
rect 0 104184 800 104304
rect 179200 103776 180000 103896
rect 0 101328 800 101448
rect 179200 101192 180000 101312
rect 0 98472 800 98592
rect 179200 98608 180000 98728
rect 179200 96024 180000 96144
rect 0 95616 800 95736
rect 179200 93440 180000 93560
rect 0 92760 800 92880
rect 179200 90856 180000 90976
rect 0 89904 800 90024
rect 179200 88272 180000 88392
rect 0 87048 800 87168
rect 179200 85688 180000 85808
rect 0 84192 800 84312
rect 179200 83104 180000 83224
rect 0 81336 800 81456
rect 179200 80520 180000 80640
rect 0 78480 800 78600
rect 179200 77936 180000 78056
rect 0 75624 800 75744
rect 179200 75352 180000 75472
rect 0 72768 800 72888
rect 179200 72768 180000 72888
rect 179200 70184 180000 70304
rect 0 69912 800 70032
rect 179200 67600 180000 67720
rect 0 67056 800 67176
rect 179200 65016 180000 65136
rect 0 64200 800 64320
rect 179200 62432 180000 62552
rect 0 61344 800 61464
rect 179200 59848 180000 59968
rect 0 58488 800 58608
rect 179200 57264 180000 57384
rect 0 55632 800 55752
rect 179200 54680 180000 54800
rect 0 52776 800 52896
rect 179200 52096 180000 52216
rect 0 49920 800 50040
rect 179200 49512 180000 49632
rect 0 47064 800 47184
rect 179200 46928 180000 47048
rect 0 44208 800 44328
rect 179200 44344 180000 44464
rect 179200 41760 180000 41880
rect 0 41352 800 41472
rect 179200 39176 180000 39296
rect 0 38496 800 38616
rect 179200 36592 180000 36712
rect 0 35640 800 35760
rect 179200 34008 180000 34128
rect 0 32784 800 32904
rect 179200 31424 180000 31544
rect 0 29928 800 30048
rect 179200 28840 180000 28960
rect 0 27072 800 27192
rect 179200 26256 180000 26376
rect 0 24216 800 24336
rect 179200 23672 180000 23792
rect 0 21360 800 21480
rect 179200 21088 180000 21208
rect 0 18504 800 18624
rect 179200 18504 180000 18624
rect 179200 15920 180000 16040
rect 0 15648 800 15768
rect 179200 13336 180000 13456
rect 0 12792 800 12912
rect 179200 10752 180000 10872
rect 0 9936 800 10056
rect 179200 8168 180000 8288
rect 0 7080 800 7200
rect 179200 5584 180000 5704
rect 0 4224 800 4344
rect 179200 3000 180000 3120
rect 0 1368 800 1488
<< obsm3 >>
rect 880 118384 179200 118557
rect 800 116896 179200 118384
rect 800 116616 179120 116896
rect 800 115808 179200 116616
rect 880 115528 179200 115808
rect 800 114312 179200 115528
rect 800 114032 179120 114312
rect 800 112952 179200 114032
rect 880 112672 179200 112952
rect 800 111728 179200 112672
rect 800 111448 179120 111728
rect 800 110096 179200 111448
rect 880 109816 179200 110096
rect 800 109144 179200 109816
rect 800 108864 179120 109144
rect 800 107240 179200 108864
rect 880 106960 179200 107240
rect 800 106560 179200 106960
rect 800 106280 179120 106560
rect 800 104384 179200 106280
rect 880 104104 179200 104384
rect 800 103976 179200 104104
rect 800 103696 179120 103976
rect 800 101528 179200 103696
rect 880 101392 179200 101528
rect 880 101248 179120 101392
rect 800 101112 179120 101248
rect 800 98808 179200 101112
rect 800 98672 179120 98808
rect 880 98528 179120 98672
rect 880 98392 179200 98528
rect 800 96224 179200 98392
rect 800 95944 179120 96224
rect 800 95816 179200 95944
rect 880 95536 179200 95816
rect 800 93640 179200 95536
rect 800 93360 179120 93640
rect 800 92960 179200 93360
rect 880 92680 179200 92960
rect 800 91056 179200 92680
rect 800 90776 179120 91056
rect 800 90104 179200 90776
rect 880 89824 179200 90104
rect 800 88472 179200 89824
rect 800 88192 179120 88472
rect 800 87248 179200 88192
rect 880 86968 179200 87248
rect 800 85888 179200 86968
rect 800 85608 179120 85888
rect 800 84392 179200 85608
rect 880 84112 179200 84392
rect 800 83304 179200 84112
rect 800 83024 179120 83304
rect 800 81536 179200 83024
rect 880 81256 179200 81536
rect 800 80720 179200 81256
rect 800 80440 179120 80720
rect 800 78680 179200 80440
rect 880 78400 179200 78680
rect 800 78136 179200 78400
rect 800 77856 179120 78136
rect 800 75824 179200 77856
rect 880 75552 179200 75824
rect 880 75544 179120 75552
rect 800 75272 179120 75544
rect 800 72968 179200 75272
rect 880 72688 179120 72968
rect 800 70384 179200 72688
rect 800 70112 179120 70384
rect 880 70104 179120 70112
rect 880 69832 179200 70104
rect 800 67800 179200 69832
rect 800 67520 179120 67800
rect 800 67256 179200 67520
rect 880 66976 179200 67256
rect 800 65216 179200 66976
rect 800 64936 179120 65216
rect 800 64400 179200 64936
rect 880 64120 179200 64400
rect 800 62632 179200 64120
rect 800 62352 179120 62632
rect 800 61544 179200 62352
rect 880 61264 179200 61544
rect 800 60048 179200 61264
rect 800 59768 179120 60048
rect 800 58688 179200 59768
rect 880 58408 179200 58688
rect 800 57464 179200 58408
rect 800 57184 179120 57464
rect 800 55832 179200 57184
rect 880 55552 179200 55832
rect 800 54880 179200 55552
rect 800 54600 179120 54880
rect 800 52976 179200 54600
rect 880 52696 179200 52976
rect 800 52296 179200 52696
rect 800 52016 179120 52296
rect 800 50120 179200 52016
rect 880 49840 179200 50120
rect 800 49712 179200 49840
rect 800 49432 179120 49712
rect 800 47264 179200 49432
rect 880 47128 179200 47264
rect 880 46984 179120 47128
rect 800 46848 179120 46984
rect 800 44544 179200 46848
rect 800 44408 179120 44544
rect 880 44264 179120 44408
rect 880 44128 179200 44264
rect 800 41960 179200 44128
rect 800 41680 179120 41960
rect 800 41552 179200 41680
rect 880 41272 179200 41552
rect 800 39376 179200 41272
rect 800 39096 179120 39376
rect 800 38696 179200 39096
rect 880 38416 179200 38696
rect 800 36792 179200 38416
rect 800 36512 179120 36792
rect 800 35840 179200 36512
rect 880 35560 179200 35840
rect 800 34208 179200 35560
rect 800 33928 179120 34208
rect 800 32984 179200 33928
rect 880 32704 179200 32984
rect 800 31624 179200 32704
rect 800 31344 179120 31624
rect 800 30128 179200 31344
rect 880 29848 179200 30128
rect 800 29040 179200 29848
rect 800 28760 179120 29040
rect 800 27272 179200 28760
rect 880 26992 179200 27272
rect 800 26456 179200 26992
rect 800 26176 179120 26456
rect 800 24416 179200 26176
rect 880 24136 179200 24416
rect 800 23872 179200 24136
rect 800 23592 179120 23872
rect 800 21560 179200 23592
rect 880 21288 179200 21560
rect 880 21280 179120 21288
rect 800 21008 179120 21280
rect 800 18704 179200 21008
rect 880 18424 179120 18704
rect 800 16120 179200 18424
rect 800 15848 179120 16120
rect 880 15840 179120 15848
rect 880 15568 179200 15840
rect 800 13536 179200 15568
rect 800 13256 179120 13536
rect 800 12992 179200 13256
rect 880 12712 179200 12992
rect 800 10952 179200 12712
rect 800 10672 179120 10952
rect 800 10136 179200 10672
rect 880 9856 179200 10136
rect 800 8368 179200 9856
rect 800 8088 179120 8368
rect 800 7280 179200 8088
rect 880 7000 179200 7280
rect 800 5784 179200 7000
rect 800 5504 179120 5784
rect 800 4424 179200 5504
rect 880 4144 179200 4424
rect 800 3200 179200 4144
rect 800 2920 179120 3200
rect 800 1568 179200 2920
rect 880 1395 179200 1568
<< metal4 >>
rect 4208 2128 4528 117552
rect 19568 2128 19888 117552
rect 34928 2128 35248 117552
rect 50288 2128 50608 117552
rect 65648 2128 65968 117552
rect 81008 2128 81328 117552
rect 96368 2128 96688 117552
rect 111728 2128 112048 117552
rect 127088 2128 127408 117552
rect 142448 2128 142768 117552
rect 157808 2128 158128 117552
rect 173168 2128 173488 117552
<< obsm4 >>
rect 48083 44779 50208 117197
rect 50688 44779 65568 117197
rect 66048 44779 80928 117197
rect 81408 44779 84029 117197
<< labels >>
rlabel metal3 s 179200 3000 180000 3120 6 io_in[0]
port 1 nsew signal input
rlabel metal3 s 179200 80520 180000 80640 6 io_in[10]
port 2 nsew signal input
rlabel metal3 s 179200 88272 180000 88392 6 io_in[11]
port 3 nsew signal input
rlabel metal3 s 179200 96024 180000 96144 6 io_in[12]
port 4 nsew signal input
rlabel metal3 s 179200 103776 180000 103896 6 io_in[13]
port 5 nsew signal input
rlabel metal3 s 179200 111528 180000 111648 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 176014 119200 176070 120000 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 156142 119200 156198 120000 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 136270 119200 136326 120000 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 116398 119200 116454 120000 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 96526 119200 96582 120000 6 io_in[19]
port 11 nsew signal input
rlabel metal3 s 179200 10752 180000 10872 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 76654 119200 76710 120000 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 56782 119200 56838 120000 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 36910 119200 36966 120000 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 17038 119200 17094 120000 6 io_in[23]
port 16 nsew signal input
rlabel metal3 s 0 118464 800 118584 6 io_in[24]
port 17 nsew signal input
rlabel metal3 s 0 109896 800 110016 6 io_in[25]
port 18 nsew signal input
rlabel metal3 s 0 101328 800 101448 6 io_in[26]
port 19 nsew signal input
rlabel metal3 s 0 92760 800 92880 6 io_in[27]
port 20 nsew signal input
rlabel metal3 s 0 84192 800 84312 6 io_in[28]
port 21 nsew signal input
rlabel metal3 s 0 75624 800 75744 6 io_in[29]
port 22 nsew signal input
rlabel metal3 s 179200 18504 180000 18624 6 io_in[2]
port 23 nsew signal input
rlabel metal3 s 0 67056 800 67176 6 io_in[30]
port 24 nsew signal input
rlabel metal3 s 0 58488 800 58608 6 io_in[31]
port 25 nsew signal input
rlabel metal3 s 0 49920 800 50040 6 io_in[32]
port 26 nsew signal input
rlabel metal3 s 0 41352 800 41472 6 io_in[33]
port 27 nsew signal input
rlabel metal3 s 0 32784 800 32904 6 io_in[34]
port 28 nsew signal input
rlabel metal3 s 0 24216 800 24336 6 io_in[35]
port 29 nsew signal input
rlabel metal3 s 0 15648 800 15768 6 io_in[36]
port 30 nsew signal input
rlabel metal3 s 0 7080 800 7200 6 io_in[37]
port 31 nsew signal input
rlabel metal3 s 179200 26256 180000 26376 6 io_in[3]
port 32 nsew signal input
rlabel metal3 s 179200 34008 180000 34128 6 io_in[4]
port 33 nsew signal input
rlabel metal3 s 179200 41760 180000 41880 6 io_in[5]
port 34 nsew signal input
rlabel metal3 s 179200 49512 180000 49632 6 io_in[6]
port 35 nsew signal input
rlabel metal3 s 179200 57264 180000 57384 6 io_in[7]
port 36 nsew signal input
rlabel metal3 s 179200 65016 180000 65136 6 io_in[8]
port 37 nsew signal input
rlabel metal3 s 179200 72768 180000 72888 6 io_in[9]
port 38 nsew signal input
rlabel metal3 s 179200 8168 180000 8288 6 io_oeb[0]
port 39 nsew signal output
rlabel metal3 s 179200 85688 180000 85808 6 io_oeb[10]
port 40 nsew signal output
rlabel metal3 s 179200 93440 180000 93560 6 io_oeb[11]
port 41 nsew signal output
rlabel metal3 s 179200 101192 180000 101312 6 io_oeb[12]
port 42 nsew signal output
rlabel metal3 s 179200 108944 180000 109064 6 io_oeb[13]
port 43 nsew signal output
rlabel metal3 s 179200 116696 180000 116816 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 162766 119200 162822 120000 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 142894 119200 142950 120000 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 123022 119200 123078 120000 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 103150 119200 103206 120000 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 83278 119200 83334 120000 6 io_oeb[19]
port 49 nsew signal output
rlabel metal3 s 179200 15920 180000 16040 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 63406 119200 63462 120000 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 43534 119200 43590 120000 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 23662 119200 23718 120000 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 3790 119200 3846 120000 6 io_oeb[23]
port 54 nsew signal output
rlabel metal3 s 0 112752 800 112872 6 io_oeb[24]
port 55 nsew signal output
rlabel metal3 s 0 104184 800 104304 6 io_oeb[25]
port 56 nsew signal output
rlabel metal3 s 0 95616 800 95736 6 io_oeb[26]
port 57 nsew signal output
rlabel metal3 s 0 87048 800 87168 6 io_oeb[27]
port 58 nsew signal output
rlabel metal3 s 0 78480 800 78600 6 io_oeb[28]
port 59 nsew signal output
rlabel metal3 s 0 69912 800 70032 6 io_oeb[29]
port 60 nsew signal output
rlabel metal3 s 179200 23672 180000 23792 6 io_oeb[2]
port 61 nsew signal output
rlabel metal3 s 0 61344 800 61464 6 io_oeb[30]
port 62 nsew signal output
rlabel metal3 s 0 52776 800 52896 6 io_oeb[31]
port 63 nsew signal output
rlabel metal3 s 0 44208 800 44328 6 io_oeb[32]
port 64 nsew signal output
rlabel metal3 s 0 35640 800 35760 6 io_oeb[33]
port 65 nsew signal output
rlabel metal3 s 0 27072 800 27192 6 io_oeb[34]
port 66 nsew signal output
rlabel metal3 s 0 18504 800 18624 6 io_oeb[35]
port 67 nsew signal output
rlabel metal3 s 0 9936 800 10056 6 io_oeb[36]
port 68 nsew signal output
rlabel metal3 s 0 1368 800 1488 6 io_oeb[37]
port 69 nsew signal output
rlabel metal3 s 179200 31424 180000 31544 6 io_oeb[3]
port 70 nsew signal output
rlabel metal3 s 179200 39176 180000 39296 6 io_oeb[4]
port 71 nsew signal output
rlabel metal3 s 179200 46928 180000 47048 6 io_oeb[5]
port 72 nsew signal output
rlabel metal3 s 179200 54680 180000 54800 6 io_oeb[6]
port 73 nsew signal output
rlabel metal3 s 179200 62432 180000 62552 6 io_oeb[7]
port 74 nsew signal output
rlabel metal3 s 179200 70184 180000 70304 6 io_oeb[8]
port 75 nsew signal output
rlabel metal3 s 179200 77936 180000 78056 6 io_oeb[9]
port 76 nsew signal output
rlabel metal3 s 179200 5584 180000 5704 6 io_out[0]
port 77 nsew signal output
rlabel metal3 s 179200 83104 180000 83224 6 io_out[10]
port 78 nsew signal output
rlabel metal3 s 179200 90856 180000 90976 6 io_out[11]
port 79 nsew signal output
rlabel metal3 s 179200 98608 180000 98728 6 io_out[12]
port 80 nsew signal output
rlabel metal3 s 179200 106360 180000 106480 6 io_out[13]
port 81 nsew signal output
rlabel metal3 s 179200 114112 180000 114232 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 169390 119200 169446 120000 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 149518 119200 149574 120000 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 129646 119200 129702 120000 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 109774 119200 109830 120000 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 89902 119200 89958 120000 6 io_out[19]
port 87 nsew signal output
rlabel metal3 s 179200 13336 180000 13456 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 70030 119200 70086 120000 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 50158 119200 50214 120000 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 30286 119200 30342 120000 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 10414 119200 10470 120000 6 io_out[23]
port 92 nsew signal output
rlabel metal3 s 0 115608 800 115728 6 io_out[24]
port 93 nsew signal output
rlabel metal3 s 0 107040 800 107160 6 io_out[25]
port 94 nsew signal output
rlabel metal3 s 0 98472 800 98592 6 io_out[26]
port 95 nsew signal output
rlabel metal3 s 0 89904 800 90024 6 io_out[27]
port 96 nsew signal output
rlabel metal3 s 0 81336 800 81456 6 io_out[28]
port 97 nsew signal output
rlabel metal3 s 0 72768 800 72888 6 io_out[29]
port 98 nsew signal output
rlabel metal3 s 179200 21088 180000 21208 6 io_out[2]
port 99 nsew signal output
rlabel metal3 s 0 64200 800 64320 6 io_out[30]
port 100 nsew signal output
rlabel metal3 s 0 55632 800 55752 6 io_out[31]
port 101 nsew signal output
rlabel metal3 s 0 47064 800 47184 6 io_out[32]
port 102 nsew signal output
rlabel metal3 s 0 38496 800 38616 6 io_out[33]
port 103 nsew signal output
rlabel metal3 s 0 29928 800 30048 6 io_out[34]
port 104 nsew signal output
rlabel metal3 s 0 21360 800 21480 6 io_out[35]
port 105 nsew signal output
rlabel metal3 s 0 12792 800 12912 6 io_out[36]
port 106 nsew signal output
rlabel metal3 s 0 4224 800 4344 6 io_out[37]
port 107 nsew signal output
rlabel metal3 s 179200 28840 180000 28960 6 io_out[3]
port 108 nsew signal output
rlabel metal3 s 179200 36592 180000 36712 6 io_out[4]
port 109 nsew signal output
rlabel metal3 s 179200 44344 180000 44464 6 io_out[5]
port 110 nsew signal output
rlabel metal3 s 179200 52096 180000 52216 6 io_out[6]
port 111 nsew signal output
rlabel metal3 s 179200 59848 180000 59968 6 io_out[7]
port 112 nsew signal output
rlabel metal3 s 179200 67600 180000 67720 6 io_out[8]
port 113 nsew signal output
rlabel metal3 s 179200 75352 180000 75472 6 io_out[9]
port 114 nsew signal output
rlabel metal2 s 65338 0 65394 800 6 la_data_in[0]
port 115 nsew signal input
rlabel metal2 s 70858 0 70914 800 6 la_data_in[10]
port 116 nsew signal input
rlabel metal2 s 71410 0 71466 800 6 la_data_in[11]
port 117 nsew signal input
rlabel metal2 s 71962 0 72018 800 6 la_data_in[12]
port 118 nsew signal input
rlabel metal2 s 72514 0 72570 800 6 la_data_in[13]
port 119 nsew signal input
rlabel metal2 s 73066 0 73122 800 6 la_data_in[14]
port 120 nsew signal input
rlabel metal2 s 73618 0 73674 800 6 la_data_in[15]
port 121 nsew signal input
rlabel metal2 s 74170 0 74226 800 6 la_data_in[16]
port 122 nsew signal input
rlabel metal2 s 74722 0 74778 800 6 la_data_in[17]
port 123 nsew signal input
rlabel metal2 s 75274 0 75330 800 6 la_data_in[18]
port 124 nsew signal input
rlabel metal2 s 75826 0 75882 800 6 la_data_in[19]
port 125 nsew signal input
rlabel metal2 s 65890 0 65946 800 6 la_data_in[1]
port 126 nsew signal input
rlabel metal2 s 76378 0 76434 800 6 la_data_in[20]
port 127 nsew signal input
rlabel metal2 s 76930 0 76986 800 6 la_data_in[21]
port 128 nsew signal input
rlabel metal2 s 77482 0 77538 800 6 la_data_in[22]
port 129 nsew signal input
rlabel metal2 s 78034 0 78090 800 6 la_data_in[23]
port 130 nsew signal input
rlabel metal2 s 78586 0 78642 800 6 la_data_in[24]
port 131 nsew signal input
rlabel metal2 s 79138 0 79194 800 6 la_data_in[25]
port 132 nsew signal input
rlabel metal2 s 79690 0 79746 800 6 la_data_in[26]
port 133 nsew signal input
rlabel metal2 s 80242 0 80298 800 6 la_data_in[27]
port 134 nsew signal input
rlabel metal2 s 80794 0 80850 800 6 la_data_in[28]
port 135 nsew signal input
rlabel metal2 s 81346 0 81402 800 6 la_data_in[29]
port 136 nsew signal input
rlabel metal2 s 66442 0 66498 800 6 la_data_in[2]
port 137 nsew signal input
rlabel metal2 s 81898 0 81954 800 6 la_data_in[30]
port 138 nsew signal input
rlabel metal2 s 82450 0 82506 800 6 la_data_in[31]
port 139 nsew signal input
rlabel metal2 s 83002 0 83058 800 6 la_data_in[32]
port 140 nsew signal input
rlabel metal2 s 83554 0 83610 800 6 la_data_in[33]
port 141 nsew signal input
rlabel metal2 s 84106 0 84162 800 6 la_data_in[34]
port 142 nsew signal input
rlabel metal2 s 84658 0 84714 800 6 la_data_in[35]
port 143 nsew signal input
rlabel metal2 s 85210 0 85266 800 6 la_data_in[36]
port 144 nsew signal input
rlabel metal2 s 85762 0 85818 800 6 la_data_in[37]
port 145 nsew signal input
rlabel metal2 s 86314 0 86370 800 6 la_data_in[38]
port 146 nsew signal input
rlabel metal2 s 86866 0 86922 800 6 la_data_in[39]
port 147 nsew signal input
rlabel metal2 s 66994 0 67050 800 6 la_data_in[3]
port 148 nsew signal input
rlabel metal2 s 87418 0 87474 800 6 la_data_in[40]
port 149 nsew signal input
rlabel metal2 s 87970 0 88026 800 6 la_data_in[41]
port 150 nsew signal input
rlabel metal2 s 88522 0 88578 800 6 la_data_in[42]
port 151 nsew signal input
rlabel metal2 s 89074 0 89130 800 6 la_data_in[43]
port 152 nsew signal input
rlabel metal2 s 89626 0 89682 800 6 la_data_in[44]
port 153 nsew signal input
rlabel metal2 s 90178 0 90234 800 6 la_data_in[45]
port 154 nsew signal input
rlabel metal2 s 90730 0 90786 800 6 la_data_in[46]
port 155 nsew signal input
rlabel metal2 s 91282 0 91338 800 6 la_data_in[47]
port 156 nsew signal input
rlabel metal2 s 91834 0 91890 800 6 la_data_in[48]
port 157 nsew signal input
rlabel metal2 s 92386 0 92442 800 6 la_data_in[49]
port 158 nsew signal input
rlabel metal2 s 67546 0 67602 800 6 la_data_in[4]
port 159 nsew signal input
rlabel metal2 s 92938 0 92994 800 6 la_data_in[50]
port 160 nsew signal input
rlabel metal2 s 93490 0 93546 800 6 la_data_in[51]
port 161 nsew signal input
rlabel metal2 s 94042 0 94098 800 6 la_data_in[52]
port 162 nsew signal input
rlabel metal2 s 94594 0 94650 800 6 la_data_in[53]
port 163 nsew signal input
rlabel metal2 s 95146 0 95202 800 6 la_data_in[54]
port 164 nsew signal input
rlabel metal2 s 95698 0 95754 800 6 la_data_in[55]
port 165 nsew signal input
rlabel metal2 s 96250 0 96306 800 6 la_data_in[56]
port 166 nsew signal input
rlabel metal2 s 96802 0 96858 800 6 la_data_in[57]
port 167 nsew signal input
rlabel metal2 s 97354 0 97410 800 6 la_data_in[58]
port 168 nsew signal input
rlabel metal2 s 97906 0 97962 800 6 la_data_in[59]
port 169 nsew signal input
rlabel metal2 s 68098 0 68154 800 6 la_data_in[5]
port 170 nsew signal input
rlabel metal2 s 98458 0 98514 800 6 la_data_in[60]
port 171 nsew signal input
rlabel metal2 s 99010 0 99066 800 6 la_data_in[61]
port 172 nsew signal input
rlabel metal2 s 99562 0 99618 800 6 la_data_in[62]
port 173 nsew signal input
rlabel metal2 s 100114 0 100170 800 6 la_data_in[63]
port 174 nsew signal input
rlabel metal2 s 68650 0 68706 800 6 la_data_in[6]
port 175 nsew signal input
rlabel metal2 s 69202 0 69258 800 6 la_data_in[7]
port 176 nsew signal input
rlabel metal2 s 69754 0 69810 800 6 la_data_in[8]
port 177 nsew signal input
rlabel metal2 s 70306 0 70362 800 6 la_data_in[9]
port 178 nsew signal input
rlabel metal2 s 100666 0 100722 800 6 la_data_out[0]
port 179 nsew signal output
rlabel metal2 s 106186 0 106242 800 6 la_data_out[10]
port 180 nsew signal output
rlabel metal2 s 106738 0 106794 800 6 la_data_out[11]
port 181 nsew signal output
rlabel metal2 s 107290 0 107346 800 6 la_data_out[12]
port 182 nsew signal output
rlabel metal2 s 107842 0 107898 800 6 la_data_out[13]
port 183 nsew signal output
rlabel metal2 s 108394 0 108450 800 6 la_data_out[14]
port 184 nsew signal output
rlabel metal2 s 108946 0 109002 800 6 la_data_out[15]
port 185 nsew signal output
rlabel metal2 s 109498 0 109554 800 6 la_data_out[16]
port 186 nsew signal output
rlabel metal2 s 110050 0 110106 800 6 la_data_out[17]
port 187 nsew signal output
rlabel metal2 s 110602 0 110658 800 6 la_data_out[18]
port 188 nsew signal output
rlabel metal2 s 111154 0 111210 800 6 la_data_out[19]
port 189 nsew signal output
rlabel metal2 s 101218 0 101274 800 6 la_data_out[1]
port 190 nsew signal output
rlabel metal2 s 111706 0 111762 800 6 la_data_out[20]
port 191 nsew signal output
rlabel metal2 s 112258 0 112314 800 6 la_data_out[21]
port 192 nsew signal output
rlabel metal2 s 112810 0 112866 800 6 la_data_out[22]
port 193 nsew signal output
rlabel metal2 s 113362 0 113418 800 6 la_data_out[23]
port 194 nsew signal output
rlabel metal2 s 113914 0 113970 800 6 la_data_out[24]
port 195 nsew signal output
rlabel metal2 s 114466 0 114522 800 6 la_data_out[25]
port 196 nsew signal output
rlabel metal2 s 115018 0 115074 800 6 la_data_out[26]
port 197 nsew signal output
rlabel metal2 s 115570 0 115626 800 6 la_data_out[27]
port 198 nsew signal output
rlabel metal2 s 116122 0 116178 800 6 la_data_out[28]
port 199 nsew signal output
rlabel metal2 s 116674 0 116730 800 6 la_data_out[29]
port 200 nsew signal output
rlabel metal2 s 101770 0 101826 800 6 la_data_out[2]
port 201 nsew signal output
rlabel metal2 s 117226 0 117282 800 6 la_data_out[30]
port 202 nsew signal output
rlabel metal2 s 117778 0 117834 800 6 la_data_out[31]
port 203 nsew signal output
rlabel metal2 s 118330 0 118386 800 6 la_data_out[32]
port 204 nsew signal output
rlabel metal2 s 118882 0 118938 800 6 la_data_out[33]
port 205 nsew signal output
rlabel metal2 s 119434 0 119490 800 6 la_data_out[34]
port 206 nsew signal output
rlabel metal2 s 119986 0 120042 800 6 la_data_out[35]
port 207 nsew signal output
rlabel metal2 s 120538 0 120594 800 6 la_data_out[36]
port 208 nsew signal output
rlabel metal2 s 121090 0 121146 800 6 la_data_out[37]
port 209 nsew signal output
rlabel metal2 s 121642 0 121698 800 6 la_data_out[38]
port 210 nsew signal output
rlabel metal2 s 122194 0 122250 800 6 la_data_out[39]
port 211 nsew signal output
rlabel metal2 s 102322 0 102378 800 6 la_data_out[3]
port 212 nsew signal output
rlabel metal2 s 122746 0 122802 800 6 la_data_out[40]
port 213 nsew signal output
rlabel metal2 s 123298 0 123354 800 6 la_data_out[41]
port 214 nsew signal output
rlabel metal2 s 123850 0 123906 800 6 la_data_out[42]
port 215 nsew signal output
rlabel metal2 s 124402 0 124458 800 6 la_data_out[43]
port 216 nsew signal output
rlabel metal2 s 124954 0 125010 800 6 la_data_out[44]
port 217 nsew signal output
rlabel metal2 s 125506 0 125562 800 6 la_data_out[45]
port 218 nsew signal output
rlabel metal2 s 126058 0 126114 800 6 la_data_out[46]
port 219 nsew signal output
rlabel metal2 s 126610 0 126666 800 6 la_data_out[47]
port 220 nsew signal output
rlabel metal2 s 127162 0 127218 800 6 la_data_out[48]
port 221 nsew signal output
rlabel metal2 s 127714 0 127770 800 6 la_data_out[49]
port 222 nsew signal output
rlabel metal2 s 102874 0 102930 800 6 la_data_out[4]
port 223 nsew signal output
rlabel metal2 s 128266 0 128322 800 6 la_data_out[50]
port 224 nsew signal output
rlabel metal2 s 128818 0 128874 800 6 la_data_out[51]
port 225 nsew signal output
rlabel metal2 s 129370 0 129426 800 6 la_data_out[52]
port 226 nsew signal output
rlabel metal2 s 129922 0 129978 800 6 la_data_out[53]
port 227 nsew signal output
rlabel metal2 s 130474 0 130530 800 6 la_data_out[54]
port 228 nsew signal output
rlabel metal2 s 131026 0 131082 800 6 la_data_out[55]
port 229 nsew signal output
rlabel metal2 s 131578 0 131634 800 6 la_data_out[56]
port 230 nsew signal output
rlabel metal2 s 132130 0 132186 800 6 la_data_out[57]
port 231 nsew signal output
rlabel metal2 s 132682 0 132738 800 6 la_data_out[58]
port 232 nsew signal output
rlabel metal2 s 133234 0 133290 800 6 la_data_out[59]
port 233 nsew signal output
rlabel metal2 s 103426 0 103482 800 6 la_data_out[5]
port 234 nsew signal output
rlabel metal2 s 133786 0 133842 800 6 la_data_out[60]
port 235 nsew signal output
rlabel metal2 s 134338 0 134394 800 6 la_data_out[61]
port 236 nsew signal output
rlabel metal2 s 134890 0 134946 800 6 la_data_out[62]
port 237 nsew signal output
rlabel metal2 s 135442 0 135498 800 6 la_data_out[63]
port 238 nsew signal output
rlabel metal2 s 103978 0 104034 800 6 la_data_out[6]
port 239 nsew signal output
rlabel metal2 s 104530 0 104586 800 6 la_data_out[7]
port 240 nsew signal output
rlabel metal2 s 105082 0 105138 800 6 la_data_out[8]
port 241 nsew signal output
rlabel metal2 s 105634 0 105690 800 6 la_data_out[9]
port 242 nsew signal output
rlabel metal2 s 135994 0 136050 800 6 la_oenb[0]
port 243 nsew signal input
rlabel metal2 s 141514 0 141570 800 6 la_oenb[10]
port 244 nsew signal input
rlabel metal2 s 142066 0 142122 800 6 la_oenb[11]
port 245 nsew signal input
rlabel metal2 s 142618 0 142674 800 6 la_oenb[12]
port 246 nsew signal input
rlabel metal2 s 143170 0 143226 800 6 la_oenb[13]
port 247 nsew signal input
rlabel metal2 s 143722 0 143778 800 6 la_oenb[14]
port 248 nsew signal input
rlabel metal2 s 144274 0 144330 800 6 la_oenb[15]
port 249 nsew signal input
rlabel metal2 s 144826 0 144882 800 6 la_oenb[16]
port 250 nsew signal input
rlabel metal2 s 145378 0 145434 800 6 la_oenb[17]
port 251 nsew signal input
rlabel metal2 s 145930 0 145986 800 6 la_oenb[18]
port 252 nsew signal input
rlabel metal2 s 146482 0 146538 800 6 la_oenb[19]
port 253 nsew signal input
rlabel metal2 s 136546 0 136602 800 6 la_oenb[1]
port 254 nsew signal input
rlabel metal2 s 147034 0 147090 800 6 la_oenb[20]
port 255 nsew signal input
rlabel metal2 s 147586 0 147642 800 6 la_oenb[21]
port 256 nsew signal input
rlabel metal2 s 148138 0 148194 800 6 la_oenb[22]
port 257 nsew signal input
rlabel metal2 s 148690 0 148746 800 6 la_oenb[23]
port 258 nsew signal input
rlabel metal2 s 149242 0 149298 800 6 la_oenb[24]
port 259 nsew signal input
rlabel metal2 s 149794 0 149850 800 6 la_oenb[25]
port 260 nsew signal input
rlabel metal2 s 150346 0 150402 800 6 la_oenb[26]
port 261 nsew signal input
rlabel metal2 s 150898 0 150954 800 6 la_oenb[27]
port 262 nsew signal input
rlabel metal2 s 151450 0 151506 800 6 la_oenb[28]
port 263 nsew signal input
rlabel metal2 s 152002 0 152058 800 6 la_oenb[29]
port 264 nsew signal input
rlabel metal2 s 137098 0 137154 800 6 la_oenb[2]
port 265 nsew signal input
rlabel metal2 s 152554 0 152610 800 6 la_oenb[30]
port 266 nsew signal input
rlabel metal2 s 153106 0 153162 800 6 la_oenb[31]
port 267 nsew signal input
rlabel metal2 s 153658 0 153714 800 6 la_oenb[32]
port 268 nsew signal input
rlabel metal2 s 154210 0 154266 800 6 la_oenb[33]
port 269 nsew signal input
rlabel metal2 s 154762 0 154818 800 6 la_oenb[34]
port 270 nsew signal input
rlabel metal2 s 155314 0 155370 800 6 la_oenb[35]
port 271 nsew signal input
rlabel metal2 s 155866 0 155922 800 6 la_oenb[36]
port 272 nsew signal input
rlabel metal2 s 156418 0 156474 800 6 la_oenb[37]
port 273 nsew signal input
rlabel metal2 s 156970 0 157026 800 6 la_oenb[38]
port 274 nsew signal input
rlabel metal2 s 157522 0 157578 800 6 la_oenb[39]
port 275 nsew signal input
rlabel metal2 s 137650 0 137706 800 6 la_oenb[3]
port 276 nsew signal input
rlabel metal2 s 158074 0 158130 800 6 la_oenb[40]
port 277 nsew signal input
rlabel metal2 s 158626 0 158682 800 6 la_oenb[41]
port 278 nsew signal input
rlabel metal2 s 159178 0 159234 800 6 la_oenb[42]
port 279 nsew signal input
rlabel metal2 s 159730 0 159786 800 6 la_oenb[43]
port 280 nsew signal input
rlabel metal2 s 160282 0 160338 800 6 la_oenb[44]
port 281 nsew signal input
rlabel metal2 s 160834 0 160890 800 6 la_oenb[45]
port 282 nsew signal input
rlabel metal2 s 161386 0 161442 800 6 la_oenb[46]
port 283 nsew signal input
rlabel metal2 s 161938 0 161994 800 6 la_oenb[47]
port 284 nsew signal input
rlabel metal2 s 162490 0 162546 800 6 la_oenb[48]
port 285 nsew signal input
rlabel metal2 s 163042 0 163098 800 6 la_oenb[49]
port 286 nsew signal input
rlabel metal2 s 138202 0 138258 800 6 la_oenb[4]
port 287 nsew signal input
rlabel metal2 s 163594 0 163650 800 6 la_oenb[50]
port 288 nsew signal input
rlabel metal2 s 164146 0 164202 800 6 la_oenb[51]
port 289 nsew signal input
rlabel metal2 s 164698 0 164754 800 6 la_oenb[52]
port 290 nsew signal input
rlabel metal2 s 165250 0 165306 800 6 la_oenb[53]
port 291 nsew signal input
rlabel metal2 s 165802 0 165858 800 6 la_oenb[54]
port 292 nsew signal input
rlabel metal2 s 166354 0 166410 800 6 la_oenb[55]
port 293 nsew signal input
rlabel metal2 s 166906 0 166962 800 6 la_oenb[56]
port 294 nsew signal input
rlabel metal2 s 167458 0 167514 800 6 la_oenb[57]
port 295 nsew signal input
rlabel metal2 s 168010 0 168066 800 6 la_oenb[58]
port 296 nsew signal input
rlabel metal2 s 168562 0 168618 800 6 la_oenb[59]
port 297 nsew signal input
rlabel metal2 s 138754 0 138810 800 6 la_oenb[5]
port 298 nsew signal input
rlabel metal2 s 169114 0 169170 800 6 la_oenb[60]
port 299 nsew signal input
rlabel metal2 s 169666 0 169722 800 6 la_oenb[61]
port 300 nsew signal input
rlabel metal2 s 170218 0 170274 800 6 la_oenb[62]
port 301 nsew signal input
rlabel metal2 s 170770 0 170826 800 6 la_oenb[63]
port 302 nsew signal input
rlabel metal2 s 139306 0 139362 800 6 la_oenb[6]
port 303 nsew signal input
rlabel metal2 s 139858 0 139914 800 6 la_oenb[7]
port 304 nsew signal input
rlabel metal2 s 140410 0 140466 800 6 la_oenb[8]
port 305 nsew signal input
rlabel metal2 s 140962 0 141018 800 6 la_oenb[9]
port 306 nsew signal input
rlabel metal2 s 171322 0 171378 800 6 user_clock2
port 307 nsew signal input
rlabel metal2 s 171874 0 171930 800 6 user_irq[0]
port 308 nsew signal output
rlabel metal2 s 172426 0 172482 800 6 user_irq[1]
port 309 nsew signal output
rlabel metal2 s 172978 0 173034 800 6 user_irq[2]
port 310 nsew signal output
rlabel metal4 s 4208 2128 4528 117552 6 vccd1
port 311 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 117552 6 vccd1
port 311 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 117552 6 vccd1
port 311 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 117552 6 vccd1
port 311 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 117552 6 vccd1
port 311 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 117552 6 vccd1
port 311 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 117552 6 vssd1
port 312 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 117552 6 vssd1
port 312 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 117552 6 vssd1
port 312 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 117552 6 vssd1
port 312 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 117552 6 vssd1
port 312 nsew ground bidirectional
rlabel metal4 s 173168 2128 173488 117552 6 vssd1
port 312 nsew ground bidirectional
rlabel metal2 s 6826 0 6882 800 6 wb_clk_i
port 313 nsew signal input
rlabel metal2 s 7378 0 7434 800 6 wb_rst_i
port 314 nsew signal input
rlabel metal2 s 7930 0 7986 800 6 wbs_ack_o
port 315 nsew signal output
rlabel metal2 s 8482 0 8538 800 6 wbs_adr_i[0]
port 316 nsew signal input
rlabel metal2 s 14002 0 14058 800 6 wbs_adr_i[10]
port 317 nsew signal input
rlabel metal2 s 14554 0 14610 800 6 wbs_adr_i[11]
port 318 nsew signal input
rlabel metal2 s 15106 0 15162 800 6 wbs_adr_i[12]
port 319 nsew signal input
rlabel metal2 s 15658 0 15714 800 6 wbs_adr_i[13]
port 320 nsew signal input
rlabel metal2 s 16210 0 16266 800 6 wbs_adr_i[14]
port 321 nsew signal input
rlabel metal2 s 16762 0 16818 800 6 wbs_adr_i[15]
port 322 nsew signal input
rlabel metal2 s 17314 0 17370 800 6 wbs_adr_i[16]
port 323 nsew signal input
rlabel metal2 s 17866 0 17922 800 6 wbs_adr_i[17]
port 324 nsew signal input
rlabel metal2 s 18418 0 18474 800 6 wbs_adr_i[18]
port 325 nsew signal input
rlabel metal2 s 18970 0 19026 800 6 wbs_adr_i[19]
port 326 nsew signal input
rlabel metal2 s 9034 0 9090 800 6 wbs_adr_i[1]
port 327 nsew signal input
rlabel metal2 s 19522 0 19578 800 6 wbs_adr_i[20]
port 328 nsew signal input
rlabel metal2 s 20074 0 20130 800 6 wbs_adr_i[21]
port 329 nsew signal input
rlabel metal2 s 20626 0 20682 800 6 wbs_adr_i[22]
port 330 nsew signal input
rlabel metal2 s 21178 0 21234 800 6 wbs_adr_i[23]
port 331 nsew signal input
rlabel metal2 s 21730 0 21786 800 6 wbs_adr_i[24]
port 332 nsew signal input
rlabel metal2 s 22282 0 22338 800 6 wbs_adr_i[25]
port 333 nsew signal input
rlabel metal2 s 22834 0 22890 800 6 wbs_adr_i[26]
port 334 nsew signal input
rlabel metal2 s 23386 0 23442 800 6 wbs_adr_i[27]
port 335 nsew signal input
rlabel metal2 s 23938 0 23994 800 6 wbs_adr_i[28]
port 336 nsew signal input
rlabel metal2 s 24490 0 24546 800 6 wbs_adr_i[29]
port 337 nsew signal input
rlabel metal2 s 9586 0 9642 800 6 wbs_adr_i[2]
port 338 nsew signal input
rlabel metal2 s 25042 0 25098 800 6 wbs_adr_i[30]
port 339 nsew signal input
rlabel metal2 s 25594 0 25650 800 6 wbs_adr_i[31]
port 340 nsew signal input
rlabel metal2 s 10138 0 10194 800 6 wbs_adr_i[3]
port 341 nsew signal input
rlabel metal2 s 10690 0 10746 800 6 wbs_adr_i[4]
port 342 nsew signal input
rlabel metal2 s 11242 0 11298 800 6 wbs_adr_i[5]
port 343 nsew signal input
rlabel metal2 s 11794 0 11850 800 6 wbs_adr_i[6]
port 344 nsew signal input
rlabel metal2 s 12346 0 12402 800 6 wbs_adr_i[7]
port 345 nsew signal input
rlabel metal2 s 12898 0 12954 800 6 wbs_adr_i[8]
port 346 nsew signal input
rlabel metal2 s 13450 0 13506 800 6 wbs_adr_i[9]
port 347 nsew signal input
rlabel metal2 s 26146 0 26202 800 6 wbs_cyc_i
port 348 nsew signal input
rlabel metal2 s 26698 0 26754 800 6 wbs_dat_i[0]
port 349 nsew signal input
rlabel metal2 s 32218 0 32274 800 6 wbs_dat_i[10]
port 350 nsew signal input
rlabel metal2 s 32770 0 32826 800 6 wbs_dat_i[11]
port 351 nsew signal input
rlabel metal2 s 33322 0 33378 800 6 wbs_dat_i[12]
port 352 nsew signal input
rlabel metal2 s 33874 0 33930 800 6 wbs_dat_i[13]
port 353 nsew signal input
rlabel metal2 s 34426 0 34482 800 6 wbs_dat_i[14]
port 354 nsew signal input
rlabel metal2 s 34978 0 35034 800 6 wbs_dat_i[15]
port 355 nsew signal input
rlabel metal2 s 35530 0 35586 800 6 wbs_dat_i[16]
port 356 nsew signal input
rlabel metal2 s 36082 0 36138 800 6 wbs_dat_i[17]
port 357 nsew signal input
rlabel metal2 s 36634 0 36690 800 6 wbs_dat_i[18]
port 358 nsew signal input
rlabel metal2 s 37186 0 37242 800 6 wbs_dat_i[19]
port 359 nsew signal input
rlabel metal2 s 27250 0 27306 800 6 wbs_dat_i[1]
port 360 nsew signal input
rlabel metal2 s 37738 0 37794 800 6 wbs_dat_i[20]
port 361 nsew signal input
rlabel metal2 s 38290 0 38346 800 6 wbs_dat_i[21]
port 362 nsew signal input
rlabel metal2 s 38842 0 38898 800 6 wbs_dat_i[22]
port 363 nsew signal input
rlabel metal2 s 39394 0 39450 800 6 wbs_dat_i[23]
port 364 nsew signal input
rlabel metal2 s 39946 0 40002 800 6 wbs_dat_i[24]
port 365 nsew signal input
rlabel metal2 s 40498 0 40554 800 6 wbs_dat_i[25]
port 366 nsew signal input
rlabel metal2 s 41050 0 41106 800 6 wbs_dat_i[26]
port 367 nsew signal input
rlabel metal2 s 41602 0 41658 800 6 wbs_dat_i[27]
port 368 nsew signal input
rlabel metal2 s 42154 0 42210 800 6 wbs_dat_i[28]
port 369 nsew signal input
rlabel metal2 s 42706 0 42762 800 6 wbs_dat_i[29]
port 370 nsew signal input
rlabel metal2 s 27802 0 27858 800 6 wbs_dat_i[2]
port 371 nsew signal input
rlabel metal2 s 43258 0 43314 800 6 wbs_dat_i[30]
port 372 nsew signal input
rlabel metal2 s 43810 0 43866 800 6 wbs_dat_i[31]
port 373 nsew signal input
rlabel metal2 s 28354 0 28410 800 6 wbs_dat_i[3]
port 374 nsew signal input
rlabel metal2 s 28906 0 28962 800 6 wbs_dat_i[4]
port 375 nsew signal input
rlabel metal2 s 29458 0 29514 800 6 wbs_dat_i[5]
port 376 nsew signal input
rlabel metal2 s 30010 0 30066 800 6 wbs_dat_i[6]
port 377 nsew signal input
rlabel metal2 s 30562 0 30618 800 6 wbs_dat_i[7]
port 378 nsew signal input
rlabel metal2 s 31114 0 31170 800 6 wbs_dat_i[8]
port 379 nsew signal input
rlabel metal2 s 31666 0 31722 800 6 wbs_dat_i[9]
port 380 nsew signal input
rlabel metal2 s 44362 0 44418 800 6 wbs_dat_o[0]
port 381 nsew signal output
rlabel metal2 s 49882 0 49938 800 6 wbs_dat_o[10]
port 382 nsew signal output
rlabel metal2 s 50434 0 50490 800 6 wbs_dat_o[11]
port 383 nsew signal output
rlabel metal2 s 50986 0 51042 800 6 wbs_dat_o[12]
port 384 nsew signal output
rlabel metal2 s 51538 0 51594 800 6 wbs_dat_o[13]
port 385 nsew signal output
rlabel metal2 s 52090 0 52146 800 6 wbs_dat_o[14]
port 386 nsew signal output
rlabel metal2 s 52642 0 52698 800 6 wbs_dat_o[15]
port 387 nsew signal output
rlabel metal2 s 53194 0 53250 800 6 wbs_dat_o[16]
port 388 nsew signal output
rlabel metal2 s 53746 0 53802 800 6 wbs_dat_o[17]
port 389 nsew signal output
rlabel metal2 s 54298 0 54354 800 6 wbs_dat_o[18]
port 390 nsew signal output
rlabel metal2 s 54850 0 54906 800 6 wbs_dat_o[19]
port 391 nsew signal output
rlabel metal2 s 44914 0 44970 800 6 wbs_dat_o[1]
port 392 nsew signal output
rlabel metal2 s 55402 0 55458 800 6 wbs_dat_o[20]
port 393 nsew signal output
rlabel metal2 s 55954 0 56010 800 6 wbs_dat_o[21]
port 394 nsew signal output
rlabel metal2 s 56506 0 56562 800 6 wbs_dat_o[22]
port 395 nsew signal output
rlabel metal2 s 57058 0 57114 800 6 wbs_dat_o[23]
port 396 nsew signal output
rlabel metal2 s 57610 0 57666 800 6 wbs_dat_o[24]
port 397 nsew signal output
rlabel metal2 s 58162 0 58218 800 6 wbs_dat_o[25]
port 398 nsew signal output
rlabel metal2 s 58714 0 58770 800 6 wbs_dat_o[26]
port 399 nsew signal output
rlabel metal2 s 59266 0 59322 800 6 wbs_dat_o[27]
port 400 nsew signal output
rlabel metal2 s 59818 0 59874 800 6 wbs_dat_o[28]
port 401 nsew signal output
rlabel metal2 s 60370 0 60426 800 6 wbs_dat_o[29]
port 402 nsew signal output
rlabel metal2 s 45466 0 45522 800 6 wbs_dat_o[2]
port 403 nsew signal output
rlabel metal2 s 60922 0 60978 800 6 wbs_dat_o[30]
port 404 nsew signal output
rlabel metal2 s 61474 0 61530 800 6 wbs_dat_o[31]
port 405 nsew signal output
rlabel metal2 s 46018 0 46074 800 6 wbs_dat_o[3]
port 406 nsew signal output
rlabel metal2 s 46570 0 46626 800 6 wbs_dat_o[4]
port 407 nsew signal output
rlabel metal2 s 47122 0 47178 800 6 wbs_dat_o[5]
port 408 nsew signal output
rlabel metal2 s 47674 0 47730 800 6 wbs_dat_o[6]
port 409 nsew signal output
rlabel metal2 s 48226 0 48282 800 6 wbs_dat_o[7]
port 410 nsew signal output
rlabel metal2 s 48778 0 48834 800 6 wbs_dat_o[8]
port 411 nsew signal output
rlabel metal2 s 49330 0 49386 800 6 wbs_dat_o[9]
port 412 nsew signal output
rlabel metal2 s 62026 0 62082 800 6 wbs_sel_i[0]
port 413 nsew signal input
rlabel metal2 s 62578 0 62634 800 6 wbs_sel_i[1]
port 414 nsew signal input
rlabel metal2 s 63130 0 63186 800 6 wbs_sel_i[2]
port 415 nsew signal input
rlabel metal2 s 63682 0 63738 800 6 wbs_sel_i[3]
port 416 nsew signal input
rlabel metal2 s 64234 0 64290 800 6 wbs_stb_i
port 417 nsew signal input
rlabel metal2 s 64786 0 64842 800 6 wbs_we_i
port 418 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 180000 120000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 15938292
string GDS_FILE /home/radhe/project/matrix_multiply_mpw8/openlane/user_proj_example/runs/22_12_18_14_28/results/signoff/user_proj_example.magic.gds
string GDS_START 774948
<< end >>

